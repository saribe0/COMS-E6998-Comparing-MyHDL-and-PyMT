//-----------------------------------------------------------------------------
// ram_0x4915ea16bef085cd
//-----------------------------------------------------------------------------
// dump-vcd: False
// verilator-xinit: zeros
`default_nettype none
module ram
(
  input  wire [   9:0] addr_a,
  input  wire [   9:0] addr_b,
  input  wire [   0:0] clk,
  input  wire [   7:0] data_a,
  input  wire [   7:0] data_b,
  output reg  [   7:0] q_a,
  output reg  [   7:0] q_b,
  input  wire [   0:0] reset,
  input  wire [   0:0] we_a,
  input  wire [   0:0] we_b
);

  // wire declarations
  wire   [   7:0] ram$000;
  wire   [   7:0] ram$001;
  wire   [   7:0] ram$002;
  wire   [   7:0] ram$003;
  wire   [   7:0] ram$004;
  wire   [   7:0] ram$005;
  wire   [   7:0] ram$006;
  wire   [   7:0] ram$007;
  wire   [   7:0] ram$008;
  wire   [   7:0] ram$009;
  wire   [   7:0] ram$010;
  wire   [   7:0] ram$011;
  wire   [   7:0] ram$012;
  wire   [   7:0] ram$013;
  wire   [   7:0] ram$014;
  wire   [   7:0] ram$015;
  wire   [   7:0] ram$016;
  wire   [   7:0] ram$017;
  wire   [   7:0] ram$018;
  wire   [   7:0] ram$019;
  wire   [   7:0] ram$020;
  wire   [   7:0] ram$021;
  wire   [   7:0] ram$022;
  wire   [   7:0] ram$023;
  wire   [   7:0] ram$024;
  wire   [   7:0] ram$025;
  wire   [   7:0] ram$026;
  wire   [   7:0] ram$027;
  wire   [   7:0] ram$028;
  wire   [   7:0] ram$029;
  wire   [   7:0] ram$030;
  wire   [   7:0] ram$031;
  wire   [   7:0] ram$032;
  wire   [   7:0] ram$033;
  wire   [   7:0] ram$034;
  wire   [   7:0] ram$035;
  wire   [   7:0] ram$036;
  wire   [   7:0] ram$037;
  wire   [   7:0] ram$038;
  wire   [   7:0] ram$039;
  wire   [   7:0] ram$040;
  wire   [   7:0] ram$041;
  wire   [   7:0] ram$042;
  wire   [   7:0] ram$043;
  wire   [   7:0] ram$044;
  wire   [   7:0] ram$045;
  wire   [   7:0] ram$046;
  wire   [   7:0] ram$047;
  wire   [   7:0] ram$048;
  wire   [   7:0] ram$049;
  wire   [   7:0] ram$050;
  wire   [   7:0] ram$051;
  wire   [   7:0] ram$052;
  wire   [   7:0] ram$053;
  wire   [   7:0] ram$054;
  wire   [   7:0] ram$055;
  wire   [   7:0] ram$056;
  wire   [   7:0] ram$057;
  wire   [   7:0] ram$058;
  wire   [   7:0] ram$059;
  wire   [   7:0] ram$060;
  wire   [   7:0] ram$061;
  wire   [   7:0] ram$062;
  wire   [   7:0] ram$063;
  wire   [   7:0] ram$064;
  wire   [   7:0] ram$065;
  wire   [   7:0] ram$066;
  wire   [   7:0] ram$067;
  wire   [   7:0] ram$068;
  wire   [   7:0] ram$069;
  wire   [   7:0] ram$070;
  wire   [   7:0] ram$071;
  wire   [   7:0] ram$072;
  wire   [   7:0] ram$073;
  wire   [   7:0] ram$074;
  wire   [   7:0] ram$075;
  wire   [   7:0] ram$076;
  wire   [   7:0] ram$077;
  wire   [   7:0] ram$078;
  wire   [   7:0] ram$079;
  wire   [   7:0] ram$080;
  wire   [   7:0] ram$081;
  wire   [   7:0] ram$082;
  wire   [   7:0] ram$083;
  wire   [   7:0] ram$084;
  wire   [   7:0] ram$085;
  wire   [   7:0] ram$086;
  wire   [   7:0] ram$087;
  wire   [   7:0] ram$088;
  wire   [   7:0] ram$089;
  wire   [   7:0] ram$090;
  wire   [   7:0] ram$091;
  wire   [   7:0] ram$092;
  wire   [   7:0] ram$093;
  wire   [   7:0] ram$094;
  wire   [   7:0] ram$095;
  wire   [   7:0] ram$096;
  wire   [   7:0] ram$097;
  wire   [   7:0] ram$098;
  wire   [   7:0] ram$099;
  wire   [   7:0] ram$100;
  wire   [   7:0] ram$101;
  wire   [   7:0] ram$102;
  wire   [   7:0] ram$103;
  wire   [   7:0] ram$104;
  wire   [   7:0] ram$105;
  wire   [   7:0] ram$106;
  wire   [   7:0] ram$107;
  wire   [   7:0] ram$108;
  wire   [   7:0] ram$109;
  wire   [   7:0] ram$110;
  wire   [   7:0] ram$111;
  wire   [   7:0] ram$112;
  wire   [   7:0] ram$113;
  wire   [   7:0] ram$114;
  wire   [   7:0] ram$115;
  wire   [   7:0] ram$116;
  wire   [   7:0] ram$117;
  wire   [   7:0] ram$118;
  wire   [   7:0] ram$119;
  wire   [   7:0] ram$120;
  wire   [   7:0] ram$121;
  wire   [   7:0] ram$122;
  wire   [   7:0] ram$123;
  wire   [   7:0] ram$124;
  wire   [   7:0] ram$125;
  wire   [   7:0] ram$126;
  wire   [   7:0] ram$127;
  wire   [   7:0] ram$128;
  wire   [   7:0] ram$129;
  wire   [   7:0] ram$130;
  wire   [   7:0] ram$131;
  wire   [   7:0] ram$132;
  wire   [   7:0] ram$133;
  wire   [   7:0] ram$134;
  wire   [   7:0] ram$135;
  wire   [   7:0] ram$136;
  wire   [   7:0] ram$137;
  wire   [   7:0] ram$138;
  wire   [   7:0] ram$139;
  wire   [   7:0] ram$140;
  wire   [   7:0] ram$141;
  wire   [   7:0] ram$142;
  wire   [   7:0] ram$143;
  wire   [   7:0] ram$144;
  wire   [   7:0] ram$145;
  wire   [   7:0] ram$146;
  wire   [   7:0] ram$147;
  wire   [   7:0] ram$148;
  wire   [   7:0] ram$149;
  wire   [   7:0] ram$150;
  wire   [   7:0] ram$151;
  wire   [   7:0] ram$152;
  wire   [   7:0] ram$153;
  wire   [   7:0] ram$154;
  wire   [   7:0] ram$155;
  wire   [   7:0] ram$156;
  wire   [   7:0] ram$157;
  wire   [   7:0] ram$158;
  wire   [   7:0] ram$159;
  wire   [   7:0] ram$160;
  wire   [   7:0] ram$161;
  wire   [   7:0] ram$162;
  wire   [   7:0] ram$163;
  wire   [   7:0] ram$164;
  wire   [   7:0] ram$165;
  wire   [   7:0] ram$166;
  wire   [   7:0] ram$167;
  wire   [   7:0] ram$168;
  wire   [   7:0] ram$169;
  wire   [   7:0] ram$170;
  wire   [   7:0] ram$171;
  wire   [   7:0] ram$172;
  wire   [   7:0] ram$173;
  wire   [   7:0] ram$174;
  wire   [   7:0] ram$175;
  wire   [   7:0] ram$176;
  wire   [   7:0] ram$177;
  wire   [   7:0] ram$178;
  wire   [   7:0] ram$179;
  wire   [   7:0] ram$180;
  wire   [   7:0] ram$181;
  wire   [   7:0] ram$182;
  wire   [   7:0] ram$183;
  wire   [   7:0] ram$184;
  wire   [   7:0] ram$185;
  wire   [   7:0] ram$186;
  wire   [   7:0] ram$187;
  wire   [   7:0] ram$188;
  wire   [   7:0] ram$189;
  wire   [   7:0] ram$190;
  wire   [   7:0] ram$191;
  wire   [   7:0] ram$192;
  wire   [   7:0] ram$193;
  wire   [   7:0] ram$194;
  wire   [   7:0] ram$195;
  wire   [   7:0] ram$196;
  wire   [   7:0] ram$197;
  wire   [   7:0] ram$198;
  wire   [   7:0] ram$199;
  wire   [   7:0] ram$200;
  wire   [   7:0] ram$201;
  wire   [   7:0] ram$202;
  wire   [   7:0] ram$203;
  wire   [   7:0] ram$204;
  wire   [   7:0] ram$205;
  wire   [   7:0] ram$206;
  wire   [   7:0] ram$207;
  wire   [   7:0] ram$208;
  wire   [   7:0] ram$209;
  wire   [   7:0] ram$210;
  wire   [   7:0] ram$211;
  wire   [   7:0] ram$212;
  wire   [   7:0] ram$213;
  wire   [   7:0] ram$214;
  wire   [   7:0] ram$215;
  wire   [   7:0] ram$216;
  wire   [   7:0] ram$217;
  wire   [   7:0] ram$218;
  wire   [   7:0] ram$219;
  wire   [   7:0] ram$220;
  wire   [   7:0] ram$221;
  wire   [   7:0] ram$222;
  wire   [   7:0] ram$223;
  wire   [   7:0] ram$224;
  wire   [   7:0] ram$225;
  wire   [   7:0] ram$226;
  wire   [   7:0] ram$227;
  wire   [   7:0] ram$228;
  wire   [   7:0] ram$229;
  wire   [   7:0] ram$230;
  wire   [   7:0] ram$231;
  wire   [   7:0] ram$232;
  wire   [   7:0] ram$233;
  wire   [   7:0] ram$234;
  wire   [   7:0] ram$235;
  wire   [   7:0] ram$236;
  wire   [   7:0] ram$237;
  wire   [   7:0] ram$238;
  wire   [   7:0] ram$239;
  wire   [   7:0] ram$240;
  wire   [   7:0] ram$241;
  wire   [   7:0] ram$242;
  wire   [   7:0] ram$243;
  wire   [   7:0] ram$244;
  wire   [   7:0] ram$245;
  wire   [   7:0] ram$246;
  wire   [   7:0] ram$247;
  wire   [   7:0] ram$248;
  wire   [   7:0] ram$249;
  wire   [   7:0] ram$250;
  wire   [   7:0] ram$251;
  wire   [   7:0] ram$252;
  wire   [   7:0] ram$253;
  wire   [   7:0] ram$254;
  wire   [   7:0] ram$255;
  wire   [   7:0] ram$256;
  wire   [   7:0] ram$257;
  wire   [   7:0] ram$258;
  wire   [   7:0] ram$259;
  wire   [   7:0] ram$260;
  wire   [   7:0] ram$261;
  wire   [   7:0] ram$262;
  wire   [   7:0] ram$263;
  wire   [   7:0] ram$264;
  wire   [   7:0] ram$265;
  wire   [   7:0] ram$266;
  wire   [   7:0] ram$267;
  wire   [   7:0] ram$268;
  wire   [   7:0] ram$269;
  wire   [   7:0] ram$270;
  wire   [   7:0] ram$271;
  wire   [   7:0] ram$272;
  wire   [   7:0] ram$273;
  wire   [   7:0] ram$274;
  wire   [   7:0] ram$275;
  wire   [   7:0] ram$276;
  wire   [   7:0] ram$277;
  wire   [   7:0] ram$278;
  wire   [   7:0] ram$279;
  wire   [   7:0] ram$280;
  wire   [   7:0] ram$281;
  wire   [   7:0] ram$282;
  wire   [   7:0] ram$283;
  wire   [   7:0] ram$284;
  wire   [   7:0] ram$285;
  wire   [   7:0] ram$286;
  wire   [   7:0] ram$287;
  wire   [   7:0] ram$288;
  wire   [   7:0] ram$289;
  wire   [   7:0] ram$290;
  wire   [   7:0] ram$291;
  wire   [   7:0] ram$292;
  wire   [   7:0] ram$293;
  wire   [   7:0] ram$294;
  wire   [   7:0] ram$295;
  wire   [   7:0] ram$296;
  wire   [   7:0] ram$297;
  wire   [   7:0] ram$298;
  wire   [   7:0] ram$299;
  wire   [   7:0] ram$300;
  wire   [   7:0] ram$301;
  wire   [   7:0] ram$302;
  wire   [   7:0] ram$303;
  wire   [   7:0] ram$304;
  wire   [   7:0] ram$305;
  wire   [   7:0] ram$306;
  wire   [   7:0] ram$307;
  wire   [   7:0] ram$308;
  wire   [   7:0] ram$309;
  wire   [   7:0] ram$310;
  wire   [   7:0] ram$311;
  wire   [   7:0] ram$312;
  wire   [   7:0] ram$313;
  wire   [   7:0] ram$314;
  wire   [   7:0] ram$315;
  wire   [   7:0] ram$316;
  wire   [   7:0] ram$317;
  wire   [   7:0] ram$318;
  wire   [   7:0] ram$319;
  wire   [   7:0] ram$320;
  wire   [   7:0] ram$321;
  wire   [   7:0] ram$322;
  wire   [   7:0] ram$323;
  wire   [   7:0] ram$324;
  wire   [   7:0] ram$325;
  wire   [   7:0] ram$326;
  wire   [   7:0] ram$327;
  wire   [   7:0] ram$328;
  wire   [   7:0] ram$329;
  wire   [   7:0] ram$330;
  wire   [   7:0] ram$331;
  wire   [   7:0] ram$332;
  wire   [   7:0] ram$333;
  wire   [   7:0] ram$334;
  wire   [   7:0] ram$335;
  wire   [   7:0] ram$336;
  wire   [   7:0] ram$337;
  wire   [   7:0] ram$338;
  wire   [   7:0] ram$339;
  wire   [   7:0] ram$340;
  wire   [   7:0] ram$341;
  wire   [   7:0] ram$342;
  wire   [   7:0] ram$343;
  wire   [   7:0] ram$344;
  wire   [   7:0] ram$345;
  wire   [   7:0] ram$346;
  wire   [   7:0] ram$347;
  wire   [   7:0] ram$348;
  wire   [   7:0] ram$349;
  wire   [   7:0] ram$350;
  wire   [   7:0] ram$351;
  wire   [   7:0] ram$352;
  wire   [   7:0] ram$353;
  wire   [   7:0] ram$354;
  wire   [   7:0] ram$355;
  wire   [   7:0] ram$356;
  wire   [   7:0] ram$357;
  wire   [   7:0] ram$358;
  wire   [   7:0] ram$359;
  wire   [   7:0] ram$360;
  wire   [   7:0] ram$361;
  wire   [   7:0] ram$362;
  wire   [   7:0] ram$363;
  wire   [   7:0] ram$364;
  wire   [   7:0] ram$365;
  wire   [   7:0] ram$366;
  wire   [   7:0] ram$367;
  wire   [   7:0] ram$368;
  wire   [   7:0] ram$369;
  wire   [   7:0] ram$370;
  wire   [   7:0] ram$371;
  wire   [   7:0] ram$372;
  wire   [   7:0] ram$373;
  wire   [   7:0] ram$374;
  wire   [   7:0] ram$375;
  wire   [   7:0] ram$376;
  wire   [   7:0] ram$377;
  wire   [   7:0] ram$378;
  wire   [   7:0] ram$379;
  wire   [   7:0] ram$380;
  wire   [   7:0] ram$381;
  wire   [   7:0] ram$382;
  wire   [   7:0] ram$383;
  wire   [   7:0] ram$384;
  wire   [   7:0] ram$385;
  wire   [   7:0] ram$386;
  wire   [   7:0] ram$387;
  wire   [   7:0] ram$388;
  wire   [   7:0] ram$389;
  wire   [   7:0] ram$390;
  wire   [   7:0] ram$391;
  wire   [   7:0] ram$392;
  wire   [   7:0] ram$393;
  wire   [   7:0] ram$394;
  wire   [   7:0] ram$395;
  wire   [   7:0] ram$396;
  wire   [   7:0] ram$397;
  wire   [   7:0] ram$398;
  wire   [   7:0] ram$399;
  wire   [   7:0] ram$400;
  wire   [   7:0] ram$401;
  wire   [   7:0] ram$402;
  wire   [   7:0] ram$403;
  wire   [   7:0] ram$404;
  wire   [   7:0] ram$405;
  wire   [   7:0] ram$406;
  wire   [   7:0] ram$407;
  wire   [   7:0] ram$408;
  wire   [   7:0] ram$409;
  wire   [   7:0] ram$410;
  wire   [   7:0] ram$411;
  wire   [   7:0] ram$412;
  wire   [   7:0] ram$413;
  wire   [   7:0] ram$414;
  wire   [   7:0] ram$415;
  wire   [   7:0] ram$416;
  wire   [   7:0] ram$417;
  wire   [   7:0] ram$418;
  wire   [   7:0] ram$419;
  wire   [   7:0] ram$420;
  wire   [   7:0] ram$421;
  wire   [   7:0] ram$422;
  wire   [   7:0] ram$423;
  wire   [   7:0] ram$424;
  wire   [   7:0] ram$425;
  wire   [   7:0] ram$426;
  wire   [   7:0] ram$427;
  wire   [   7:0] ram$428;
  wire   [   7:0] ram$429;
  wire   [   7:0] ram$430;
  wire   [   7:0] ram$431;
  wire   [   7:0] ram$432;
  wire   [   7:0] ram$433;
  wire   [   7:0] ram$434;
  wire   [   7:0] ram$435;
  wire   [   7:0] ram$436;
  wire   [   7:0] ram$437;
  wire   [   7:0] ram$438;
  wire   [   7:0] ram$439;
  wire   [   7:0] ram$440;
  wire   [   7:0] ram$441;
  wire   [   7:0] ram$442;
  wire   [   7:0] ram$443;
  wire   [   7:0] ram$444;
  wire   [   7:0] ram$445;
  wire   [   7:0] ram$446;
  wire   [   7:0] ram$447;
  wire   [   7:0] ram$448;
  wire   [   7:0] ram$449;
  wire   [   7:0] ram$450;
  wire   [   7:0] ram$451;
  wire   [   7:0] ram$452;
  wire   [   7:0] ram$453;
  wire   [   7:0] ram$454;
  wire   [   7:0] ram$455;
  wire   [   7:0] ram$456;
  wire   [   7:0] ram$457;
  wire   [   7:0] ram$458;
  wire   [   7:0] ram$459;
  wire   [   7:0] ram$460;
  wire   [   7:0] ram$461;
  wire   [   7:0] ram$462;
  wire   [   7:0] ram$463;
  wire   [   7:0] ram$464;
  wire   [   7:0] ram$465;
  wire   [   7:0] ram$466;
  wire   [   7:0] ram$467;
  wire   [   7:0] ram$468;
  wire   [   7:0] ram$469;
  wire   [   7:0] ram$470;
  wire   [   7:0] ram$471;
  wire   [   7:0] ram$472;
  wire   [   7:0] ram$473;
  wire   [   7:0] ram$474;
  wire   [   7:0] ram$475;
  wire   [   7:0] ram$476;
  wire   [   7:0] ram$477;
  wire   [   7:0] ram$478;
  wire   [   7:0] ram$479;
  wire   [   7:0] ram$480;
  wire   [   7:0] ram$481;
  wire   [   7:0] ram$482;
  wire   [   7:0] ram$483;
  wire   [   7:0] ram$484;
  wire   [   7:0] ram$485;
  wire   [   7:0] ram$486;
  wire   [   7:0] ram$487;
  wire   [   7:0] ram$488;
  wire   [   7:0] ram$489;
  wire   [   7:0] ram$490;
  wire   [   7:0] ram$491;
  wire   [   7:0] ram$492;
  wire   [   7:0] ram$493;
  wire   [   7:0] ram$494;
  wire   [   7:0] ram$495;
  wire   [   7:0] ram$496;
  wire   [   7:0] ram$497;
  wire   [   7:0] ram$498;
  wire   [   7:0] ram$499;
  wire   [   7:0] ram$500;
  wire   [   7:0] ram$501;
  wire   [   7:0] ram$502;
  wire   [   7:0] ram$503;
  wire   [   7:0] ram$504;
  wire   [   7:0] ram$505;
  wire   [   7:0] ram$506;
  wire   [   7:0] ram$507;
  wire   [   7:0] ram$508;
  wire   [   7:0] ram$509;
  wire   [   7:0] ram$510;
  wire   [   7:0] ram$511;
  wire   [   7:0] ram$512;
  wire   [   7:0] ram$513;
  wire   [   7:0] ram$514;
  wire   [   7:0] ram$515;
  wire   [   7:0] ram$516;
  wire   [   7:0] ram$517;
  wire   [   7:0] ram$518;
  wire   [   7:0] ram$519;
  wire   [   7:0] ram$520;
  wire   [   7:0] ram$521;
  wire   [   7:0] ram$522;
  wire   [   7:0] ram$523;
  wire   [   7:0] ram$524;
  wire   [   7:0] ram$525;
  wire   [   7:0] ram$526;
  wire   [   7:0] ram$527;
  wire   [   7:0] ram$528;
  wire   [   7:0] ram$529;
  wire   [   7:0] ram$530;
  wire   [   7:0] ram$531;
  wire   [   7:0] ram$532;
  wire   [   7:0] ram$533;
  wire   [   7:0] ram$534;
  wire   [   7:0] ram$535;
  wire   [   7:0] ram$536;
  wire   [   7:0] ram$537;
  wire   [   7:0] ram$538;
  wire   [   7:0] ram$539;
  wire   [   7:0] ram$540;
  wire   [   7:0] ram$541;
  wire   [   7:0] ram$542;
  wire   [   7:0] ram$543;
  wire   [   7:0] ram$544;
  wire   [   7:0] ram$545;
  wire   [   7:0] ram$546;
  wire   [   7:0] ram$547;
  wire   [   7:0] ram$548;
  wire   [   7:0] ram$549;
  wire   [   7:0] ram$550;
  wire   [   7:0] ram$551;
  wire   [   7:0] ram$552;
  wire   [   7:0] ram$553;
  wire   [   7:0] ram$554;
  wire   [   7:0] ram$555;
  wire   [   7:0] ram$556;
  wire   [   7:0] ram$557;
  wire   [   7:0] ram$558;
  wire   [   7:0] ram$559;
  wire   [   7:0] ram$560;
  wire   [   7:0] ram$561;
  wire   [   7:0] ram$562;
  wire   [   7:0] ram$563;
  wire   [   7:0] ram$564;
  wire   [   7:0] ram$565;
  wire   [   7:0] ram$566;
  wire   [   7:0] ram$567;
  wire   [   7:0] ram$568;
  wire   [   7:0] ram$569;
  wire   [   7:0] ram$570;
  wire   [   7:0] ram$571;
  wire   [   7:0] ram$572;
  wire   [   7:0] ram$573;
  wire   [   7:0] ram$574;
  wire   [   7:0] ram$575;
  wire   [   7:0] ram$576;
  wire   [   7:0] ram$577;
  wire   [   7:0] ram$578;
  wire   [   7:0] ram$579;
  wire   [   7:0] ram$580;
  wire   [   7:0] ram$581;
  wire   [   7:0] ram$582;
  wire   [   7:0] ram$583;
  wire   [   7:0] ram$584;
  wire   [   7:0] ram$585;
  wire   [   7:0] ram$586;
  wire   [   7:0] ram$587;
  wire   [   7:0] ram$588;
  wire   [   7:0] ram$589;
  wire   [   7:0] ram$590;
  wire   [   7:0] ram$591;
  wire   [   7:0] ram$592;
  wire   [   7:0] ram$593;
  wire   [   7:0] ram$594;
  wire   [   7:0] ram$595;
  wire   [   7:0] ram$596;
  wire   [   7:0] ram$597;
  wire   [   7:0] ram$598;
  wire   [   7:0] ram$599;
  wire   [   7:0] ram$600;
  wire   [   7:0] ram$601;
  wire   [   7:0] ram$602;
  wire   [   7:0] ram$603;
  wire   [   7:0] ram$604;
  wire   [   7:0] ram$605;
  wire   [   7:0] ram$606;
  wire   [   7:0] ram$607;
  wire   [   7:0] ram$608;
  wire   [   7:0] ram$609;
  wire   [   7:0] ram$610;
  wire   [   7:0] ram$611;
  wire   [   7:0] ram$612;
  wire   [   7:0] ram$613;
  wire   [   7:0] ram$614;
  wire   [   7:0] ram$615;
  wire   [   7:0] ram$616;
  wire   [   7:0] ram$617;
  wire   [   7:0] ram$618;
  wire   [   7:0] ram$619;
  wire   [   7:0] ram$620;
  wire   [   7:0] ram$621;
  wire   [   7:0] ram$622;
  wire   [   7:0] ram$623;
  wire   [   7:0] ram$624;
  wire   [   7:0] ram$625;
  wire   [   7:0] ram$626;
  wire   [   7:0] ram$627;
  wire   [   7:0] ram$628;
  wire   [   7:0] ram$629;
  wire   [   7:0] ram$630;
  wire   [   7:0] ram$631;
  wire   [   7:0] ram$632;
  wire   [   7:0] ram$633;
  wire   [   7:0] ram$634;
  wire   [   7:0] ram$635;
  wire   [   7:0] ram$636;
  wire   [   7:0] ram$637;
  wire   [   7:0] ram$638;
  wire   [   7:0] ram$639;
  wire   [   7:0] ram$640;
  wire   [   7:0] ram$641;
  wire   [   7:0] ram$642;
  wire   [   7:0] ram$643;
  wire   [   7:0] ram$644;
  wire   [   7:0] ram$645;
  wire   [   7:0] ram$646;
  wire   [   7:0] ram$647;
  wire   [   7:0] ram$648;
  wire   [   7:0] ram$649;
  wire   [   7:0] ram$650;
  wire   [   7:0] ram$651;
  wire   [   7:0] ram$652;
  wire   [   7:0] ram$653;
  wire   [   7:0] ram$654;
  wire   [   7:0] ram$655;
  wire   [   7:0] ram$656;
  wire   [   7:0] ram$657;
  wire   [   7:0] ram$658;
  wire   [   7:0] ram$659;
  wire   [   7:0] ram$660;
  wire   [   7:0] ram$661;
  wire   [   7:0] ram$662;
  wire   [   7:0] ram$663;
  wire   [   7:0] ram$664;
  wire   [   7:0] ram$665;
  wire   [   7:0] ram$666;
  wire   [   7:0] ram$667;
  wire   [   7:0] ram$668;
  wire   [   7:0] ram$669;
  wire   [   7:0] ram$670;
  wire   [   7:0] ram$671;
  wire   [   7:0] ram$672;
  wire   [   7:0] ram$673;
  wire   [   7:0] ram$674;
  wire   [   7:0] ram$675;
  wire   [   7:0] ram$676;
  wire   [   7:0] ram$677;
  wire   [   7:0] ram$678;
  wire   [   7:0] ram$679;
  wire   [   7:0] ram$680;
  wire   [   7:0] ram$681;
  wire   [   7:0] ram$682;
  wire   [   7:0] ram$683;
  wire   [   7:0] ram$684;
  wire   [   7:0] ram$685;
  wire   [   7:0] ram$686;
  wire   [   7:0] ram$687;
  wire   [   7:0] ram$688;
  wire   [   7:0] ram$689;
  wire   [   7:0] ram$690;
  wire   [   7:0] ram$691;
  wire   [   7:0] ram$692;
  wire   [   7:0] ram$693;
  wire   [   7:0] ram$694;
  wire   [   7:0] ram$695;
  wire   [   7:0] ram$696;
  wire   [   7:0] ram$697;
  wire   [   7:0] ram$698;
  wire   [   7:0] ram$699;
  wire   [   7:0] ram$700;
  wire   [   7:0] ram$701;
  wire   [   7:0] ram$702;
  wire   [   7:0] ram$703;
  wire   [   7:0] ram$704;
  wire   [   7:0] ram$705;
  wire   [   7:0] ram$706;
  wire   [   7:0] ram$707;
  wire   [   7:0] ram$708;
  wire   [   7:0] ram$709;
  wire   [   7:0] ram$710;
  wire   [   7:0] ram$711;
  wire   [   7:0] ram$712;
  wire   [   7:0] ram$713;
  wire   [   7:0] ram$714;
  wire   [   7:0] ram$715;
  wire   [   7:0] ram$716;
  wire   [   7:0] ram$717;
  wire   [   7:0] ram$718;
  wire   [   7:0] ram$719;
  wire   [   7:0] ram$720;
  wire   [   7:0] ram$721;
  wire   [   7:0] ram$722;
  wire   [   7:0] ram$723;
  wire   [   7:0] ram$724;
  wire   [   7:0] ram$725;
  wire   [   7:0] ram$726;
  wire   [   7:0] ram$727;
  wire   [   7:0] ram$728;
  wire   [   7:0] ram$729;
  wire   [   7:0] ram$730;
  wire   [   7:0] ram$731;
  wire   [   7:0] ram$732;
  wire   [   7:0] ram$733;
  wire   [   7:0] ram$734;
  wire   [   7:0] ram$735;
  wire   [   7:0] ram$736;
  wire   [   7:0] ram$737;
  wire   [   7:0] ram$738;
  wire   [   7:0] ram$739;
  wire   [   7:0] ram$740;
  wire   [   7:0] ram$741;
  wire   [   7:0] ram$742;
  wire   [   7:0] ram$743;
  wire   [   7:0] ram$744;
  wire   [   7:0] ram$745;
  wire   [   7:0] ram$746;
  wire   [   7:0] ram$747;
  wire   [   7:0] ram$748;
  wire   [   7:0] ram$749;
  wire   [   7:0] ram$750;
  wire   [   7:0] ram$751;
  wire   [   7:0] ram$752;
  wire   [   7:0] ram$753;
  wire   [   7:0] ram$754;
  wire   [   7:0] ram$755;
  wire   [   7:0] ram$756;
  wire   [   7:0] ram$757;
  wire   [   7:0] ram$758;
  wire   [   7:0] ram$759;
  wire   [   7:0] ram$760;
  wire   [   7:0] ram$761;
  wire   [   7:0] ram$762;
  wire   [   7:0] ram$763;
  wire   [   7:0] ram$764;
  wire   [   7:0] ram$765;
  wire   [   7:0] ram$766;
  wire   [   7:0] ram$767;
  wire   [   7:0] ram$768;
  wire   [   7:0] ram$769;
  wire   [   7:0] ram$770;
  wire   [   7:0] ram$771;
  wire   [   7:0] ram$772;
  wire   [   7:0] ram$773;
  wire   [   7:0] ram$774;
  wire   [   7:0] ram$775;
  wire   [   7:0] ram$776;
  wire   [   7:0] ram$777;
  wire   [   7:0] ram$778;
  wire   [   7:0] ram$779;
  wire   [   7:0] ram$780;
  wire   [   7:0] ram$781;
  wire   [   7:0] ram$782;
  wire   [   7:0] ram$783;
  wire   [   7:0] ram$784;
  wire   [   7:0] ram$785;
  wire   [   7:0] ram$786;
  wire   [   7:0] ram$787;
  wire   [   7:0] ram$788;
  wire   [   7:0] ram$789;
  wire   [   7:0] ram$790;
  wire   [   7:0] ram$791;
  wire   [   7:0] ram$792;
  wire   [   7:0] ram$793;
  wire   [   7:0] ram$794;
  wire   [   7:0] ram$795;
  wire   [   7:0] ram$796;
  wire   [   7:0] ram$797;
  wire   [   7:0] ram$798;
  wire   [   7:0] ram$799;
  wire   [   7:0] ram$800;
  wire   [   7:0] ram$801;
  wire   [   7:0] ram$802;
  wire   [   7:0] ram$803;
  wire   [   7:0] ram$804;
  wire   [   7:0] ram$805;
  wire   [   7:0] ram$806;
  wire   [   7:0] ram$807;
  wire   [   7:0] ram$808;
  wire   [   7:0] ram$809;
  wire   [   7:0] ram$810;
  wire   [   7:0] ram$811;
  wire   [   7:0] ram$812;
  wire   [   7:0] ram$813;
  wire   [   7:0] ram$814;
  wire   [   7:0] ram$815;
  wire   [   7:0] ram$816;
  wire   [   7:0] ram$817;
  wire   [   7:0] ram$818;
  wire   [   7:0] ram$819;
  wire   [   7:0] ram$820;
  wire   [   7:0] ram$821;
  wire   [   7:0] ram$822;
  wire   [   7:0] ram$823;
  wire   [   7:0] ram$824;
  wire   [   7:0] ram$825;
  wire   [   7:0] ram$826;
  wire   [   7:0] ram$827;
  wire   [   7:0] ram$828;
  wire   [   7:0] ram$829;
  wire   [   7:0] ram$830;
  wire   [   7:0] ram$831;
  wire   [   7:0] ram$832;
  wire   [   7:0] ram$833;
  wire   [   7:0] ram$834;
  wire   [   7:0] ram$835;
  wire   [   7:0] ram$836;
  wire   [   7:0] ram$837;
  wire   [   7:0] ram$838;
  wire   [   7:0] ram$839;
  wire   [   7:0] ram$840;
  wire   [   7:0] ram$841;
  wire   [   7:0] ram$842;
  wire   [   7:0] ram$843;
  wire   [   7:0] ram$844;
  wire   [   7:0] ram$845;
  wire   [   7:0] ram$846;
  wire   [   7:0] ram$847;
  wire   [   7:0] ram$848;
  wire   [   7:0] ram$849;
  wire   [   7:0] ram$850;
  wire   [   7:0] ram$851;
  wire   [   7:0] ram$852;
  wire   [   7:0] ram$853;
  wire   [   7:0] ram$854;
  wire   [   7:0] ram$855;
  wire   [   7:0] ram$856;
  wire   [   7:0] ram$857;
  wire   [   7:0] ram$858;
  wire   [   7:0] ram$859;
  wire   [   7:0] ram$860;
  wire   [   7:0] ram$861;
  wire   [   7:0] ram$862;
  wire   [   7:0] ram$863;
  wire   [   7:0] ram$864;
  wire   [   7:0] ram$865;
  wire   [   7:0] ram$866;
  wire   [   7:0] ram$867;
  wire   [   7:0] ram$868;
  wire   [   7:0] ram$869;
  wire   [   7:0] ram$870;
  wire   [   7:0] ram$871;
  wire   [   7:0] ram$872;
  wire   [   7:0] ram$873;
  wire   [   7:0] ram$874;
  wire   [   7:0] ram$875;
  wire   [   7:0] ram$876;
  wire   [   7:0] ram$877;
  wire   [   7:0] ram$878;
  wire   [   7:0] ram$879;
  wire   [   7:0] ram$880;
  wire   [   7:0] ram$881;
  wire   [   7:0] ram$882;
  wire   [   7:0] ram$883;
  wire   [   7:0] ram$884;
  wire   [   7:0] ram$885;
  wire   [   7:0] ram$886;
  wire   [   7:0] ram$887;
  wire   [   7:0] ram$888;
  wire   [   7:0] ram$889;
  wire   [   7:0] ram$890;
  wire   [   7:0] ram$891;
  wire   [   7:0] ram$892;
  wire   [   7:0] ram$893;
  wire   [   7:0] ram$894;
  wire   [   7:0] ram$895;
  wire   [   7:0] ram$896;
  wire   [   7:0] ram$897;
  wire   [   7:0] ram$898;
  wire   [   7:0] ram$899;
  wire   [   7:0] ram$900;
  wire   [   7:0] ram$901;
  wire   [   7:0] ram$902;
  wire   [   7:0] ram$903;
  wire   [   7:0] ram$904;
  wire   [   7:0] ram$905;
  wire   [   7:0] ram$906;
  wire   [   7:0] ram$907;
  wire   [   7:0] ram$908;
  wire   [   7:0] ram$909;
  wire   [   7:0] ram$910;
  wire   [   7:0] ram$911;
  wire   [   7:0] ram$912;
  wire   [   7:0] ram$913;
  wire   [   7:0] ram$914;
  wire   [   7:0] ram$915;
  wire   [   7:0] ram$916;
  wire   [   7:0] ram$917;
  wire   [   7:0] ram$918;
  wire   [   7:0] ram$919;
  wire   [   7:0] ram$920;
  wire   [   7:0] ram$921;
  wire   [   7:0] ram$922;
  wire   [   7:0] ram$923;
  wire   [   7:0] ram$924;
  wire   [   7:0] ram$925;
  wire   [   7:0] ram$926;
  wire   [   7:0] ram$927;
  wire   [   7:0] ram$928;
  wire   [   7:0] ram$929;
  wire   [   7:0] ram$930;
  wire   [   7:0] ram$931;
  wire   [   7:0] ram$932;
  wire   [   7:0] ram$933;
  wire   [   7:0] ram$934;
  wire   [   7:0] ram$935;
  wire   [   7:0] ram$936;
  wire   [   7:0] ram$937;
  wire   [   7:0] ram$938;
  wire   [   7:0] ram$939;
  wire   [   7:0] ram$940;
  wire   [   7:0] ram$941;
  wire   [   7:0] ram$942;
  wire   [   7:0] ram$943;
  wire   [   7:0] ram$944;
  wire   [   7:0] ram$945;
  wire   [   7:0] ram$946;
  wire   [   7:0] ram$947;
  wire   [   7:0] ram$948;
  wire   [   7:0] ram$949;
  wire   [   7:0] ram$950;
  wire   [   7:0] ram$951;
  wire   [   7:0] ram$952;
  wire   [   7:0] ram$953;
  wire   [   7:0] ram$954;
  wire   [   7:0] ram$955;
  wire   [   7:0] ram$956;
  wire   [   7:0] ram$957;
  wire   [   7:0] ram$958;
  wire   [   7:0] ram$959;
  wire   [   7:0] ram$960;
  wire   [   7:0] ram$961;
  wire   [   7:0] ram$962;
  wire   [   7:0] ram$963;
  wire   [   7:0] ram$964;
  wire   [   7:0] ram$965;
  wire   [   7:0] ram$966;
  wire   [   7:0] ram$967;
  wire   [   7:0] ram$968;
  wire   [   7:0] ram$969;
  wire   [   7:0] ram$970;
  wire   [   7:0] ram$971;
  wire   [   7:0] ram$972;
  wire   [   7:0] ram$973;
  wire   [   7:0] ram$974;
  wire   [   7:0] ram$975;
  wire   [   7:0] ram$976;
  wire   [   7:0] ram$977;
  wire   [   7:0] ram$978;
  wire   [   7:0] ram$979;
  wire   [   7:0] ram$980;
  wire   [   7:0] ram$981;
  wire   [   7:0] ram$982;
  wire   [   7:0] ram$983;
  wire   [   7:0] ram$984;
  wire   [   7:0] ram$985;
  wire   [   7:0] ram$986;
  wire   [   7:0] ram$987;
  wire   [   7:0] ram$988;
  wire   [   7:0] ram$989;
  wire   [   7:0] ram$990;
  wire   [   7:0] ram$991;
  wire   [   7:0] ram$992;
  wire   [   7:0] ram$993;
  wire   [   7:0] ram$994;
  wire   [   7:0] ram$995;
  wire   [   7:0] ram$996;
  wire   [   7:0] ram$997;
  wire   [   7:0] ram$998;
  wire   [   7:0] ram$999;
  wire   [   7:0] ram$1000;
  wire   [   7:0] ram$1001;
  wire   [   7:0] ram$1002;
  wire   [   7:0] ram$1003;
  wire   [   7:0] ram$1004;
  wire   [   7:0] ram$1005;
  wire   [   7:0] ram$1006;
  wire   [   7:0] ram$1007;
  wire   [   7:0] ram$1008;
  wire   [   7:0] ram$1009;
  wire   [   7:0] ram$1010;
  wire   [   7:0] ram$1011;
  wire   [   7:0] ram$1012;
  wire   [   7:0] ram$1013;
  wire   [   7:0] ram$1014;
  wire   [   7:0] ram$1015;
  wire   [   7:0] ram$1016;
  wire   [   7:0] ram$1017;
  wire   [   7:0] ram$1018;
  wire   [   7:0] ram$1019;
  wire   [   7:0] ram$1020;
  wire   [   7:0] ram$1021;
  wire   [   7:0] ram$1022;
  wire   [   7:0] ram$1023;



  // array declarations
  reg    [   7:0] ram[0:1023];
  assign ram$000 = ram[  0];
  assign ram$001 = ram[  1];
  assign ram$002 = ram[  2];
  assign ram$003 = ram[  3];
  assign ram$004 = ram[  4];
  assign ram$005 = ram[  5];
  assign ram$006 = ram[  6];
  assign ram$007 = ram[  7];
  assign ram$008 = ram[  8];
  assign ram$009 = ram[  9];
  assign ram$010 = ram[ 10];
  assign ram$011 = ram[ 11];
  assign ram$012 = ram[ 12];
  assign ram$013 = ram[ 13];
  assign ram$014 = ram[ 14];
  assign ram$015 = ram[ 15];
  assign ram$016 = ram[ 16];
  assign ram$017 = ram[ 17];
  assign ram$018 = ram[ 18];
  assign ram$019 = ram[ 19];
  assign ram$020 = ram[ 20];
  assign ram$021 = ram[ 21];
  assign ram$022 = ram[ 22];
  assign ram$023 = ram[ 23];
  assign ram$024 = ram[ 24];
  assign ram$025 = ram[ 25];
  assign ram$026 = ram[ 26];
  assign ram$027 = ram[ 27];
  assign ram$028 = ram[ 28];
  assign ram$029 = ram[ 29];
  assign ram$030 = ram[ 30];
  assign ram$031 = ram[ 31];
  assign ram$032 = ram[ 32];
  assign ram$033 = ram[ 33];
  assign ram$034 = ram[ 34];
  assign ram$035 = ram[ 35];
  assign ram$036 = ram[ 36];
  assign ram$037 = ram[ 37];
  assign ram$038 = ram[ 38];
  assign ram$039 = ram[ 39];
  assign ram$040 = ram[ 40];
  assign ram$041 = ram[ 41];
  assign ram$042 = ram[ 42];
  assign ram$043 = ram[ 43];
  assign ram$044 = ram[ 44];
  assign ram$045 = ram[ 45];
  assign ram$046 = ram[ 46];
  assign ram$047 = ram[ 47];
  assign ram$048 = ram[ 48];
  assign ram$049 = ram[ 49];
  assign ram$050 = ram[ 50];
  assign ram$051 = ram[ 51];
  assign ram$052 = ram[ 52];
  assign ram$053 = ram[ 53];
  assign ram$054 = ram[ 54];
  assign ram$055 = ram[ 55];
  assign ram$056 = ram[ 56];
  assign ram$057 = ram[ 57];
  assign ram$058 = ram[ 58];
  assign ram$059 = ram[ 59];
  assign ram$060 = ram[ 60];
  assign ram$061 = ram[ 61];
  assign ram$062 = ram[ 62];
  assign ram$063 = ram[ 63];
  assign ram$064 = ram[ 64];
  assign ram$065 = ram[ 65];
  assign ram$066 = ram[ 66];
  assign ram$067 = ram[ 67];
  assign ram$068 = ram[ 68];
  assign ram$069 = ram[ 69];
  assign ram$070 = ram[ 70];
  assign ram$071 = ram[ 71];
  assign ram$072 = ram[ 72];
  assign ram$073 = ram[ 73];
  assign ram$074 = ram[ 74];
  assign ram$075 = ram[ 75];
  assign ram$076 = ram[ 76];
  assign ram$077 = ram[ 77];
  assign ram$078 = ram[ 78];
  assign ram$079 = ram[ 79];
  assign ram$080 = ram[ 80];
  assign ram$081 = ram[ 81];
  assign ram$082 = ram[ 82];
  assign ram$083 = ram[ 83];
  assign ram$084 = ram[ 84];
  assign ram$085 = ram[ 85];
  assign ram$086 = ram[ 86];
  assign ram$087 = ram[ 87];
  assign ram$088 = ram[ 88];
  assign ram$089 = ram[ 89];
  assign ram$090 = ram[ 90];
  assign ram$091 = ram[ 91];
  assign ram$092 = ram[ 92];
  assign ram$093 = ram[ 93];
  assign ram$094 = ram[ 94];
  assign ram$095 = ram[ 95];
  assign ram$096 = ram[ 96];
  assign ram$097 = ram[ 97];
  assign ram$098 = ram[ 98];
  assign ram$099 = ram[ 99];
  assign ram$100 = ram[100];
  assign ram$101 = ram[101];
  assign ram$102 = ram[102];
  assign ram$103 = ram[103];
  assign ram$104 = ram[104];
  assign ram$105 = ram[105];
  assign ram$106 = ram[106];
  assign ram$107 = ram[107];
  assign ram$108 = ram[108];
  assign ram$109 = ram[109];
  assign ram$110 = ram[110];
  assign ram$111 = ram[111];
  assign ram$112 = ram[112];
  assign ram$113 = ram[113];
  assign ram$114 = ram[114];
  assign ram$115 = ram[115];
  assign ram$116 = ram[116];
  assign ram$117 = ram[117];
  assign ram$118 = ram[118];
  assign ram$119 = ram[119];
  assign ram$120 = ram[120];
  assign ram$121 = ram[121];
  assign ram$122 = ram[122];
  assign ram$123 = ram[123];
  assign ram$124 = ram[124];
  assign ram$125 = ram[125];
  assign ram$126 = ram[126];
  assign ram$127 = ram[127];
  assign ram$128 = ram[128];
  assign ram$129 = ram[129];
  assign ram$130 = ram[130];
  assign ram$131 = ram[131];
  assign ram$132 = ram[132];
  assign ram$133 = ram[133];
  assign ram$134 = ram[134];
  assign ram$135 = ram[135];
  assign ram$136 = ram[136];
  assign ram$137 = ram[137];
  assign ram$138 = ram[138];
  assign ram$139 = ram[139];
  assign ram$140 = ram[140];
  assign ram$141 = ram[141];
  assign ram$142 = ram[142];
  assign ram$143 = ram[143];
  assign ram$144 = ram[144];
  assign ram$145 = ram[145];
  assign ram$146 = ram[146];
  assign ram$147 = ram[147];
  assign ram$148 = ram[148];
  assign ram$149 = ram[149];
  assign ram$150 = ram[150];
  assign ram$151 = ram[151];
  assign ram$152 = ram[152];
  assign ram$153 = ram[153];
  assign ram$154 = ram[154];
  assign ram$155 = ram[155];
  assign ram$156 = ram[156];
  assign ram$157 = ram[157];
  assign ram$158 = ram[158];
  assign ram$159 = ram[159];
  assign ram$160 = ram[160];
  assign ram$161 = ram[161];
  assign ram$162 = ram[162];
  assign ram$163 = ram[163];
  assign ram$164 = ram[164];
  assign ram$165 = ram[165];
  assign ram$166 = ram[166];
  assign ram$167 = ram[167];
  assign ram$168 = ram[168];
  assign ram$169 = ram[169];
  assign ram$170 = ram[170];
  assign ram$171 = ram[171];
  assign ram$172 = ram[172];
  assign ram$173 = ram[173];
  assign ram$174 = ram[174];
  assign ram$175 = ram[175];
  assign ram$176 = ram[176];
  assign ram$177 = ram[177];
  assign ram$178 = ram[178];
  assign ram$179 = ram[179];
  assign ram$180 = ram[180];
  assign ram$181 = ram[181];
  assign ram$182 = ram[182];
  assign ram$183 = ram[183];
  assign ram$184 = ram[184];
  assign ram$185 = ram[185];
  assign ram$186 = ram[186];
  assign ram$187 = ram[187];
  assign ram$188 = ram[188];
  assign ram$189 = ram[189];
  assign ram$190 = ram[190];
  assign ram$191 = ram[191];
  assign ram$192 = ram[192];
  assign ram$193 = ram[193];
  assign ram$194 = ram[194];
  assign ram$195 = ram[195];
  assign ram$196 = ram[196];
  assign ram$197 = ram[197];
  assign ram$198 = ram[198];
  assign ram$199 = ram[199];
  assign ram$200 = ram[200];
  assign ram$201 = ram[201];
  assign ram$202 = ram[202];
  assign ram$203 = ram[203];
  assign ram$204 = ram[204];
  assign ram$205 = ram[205];
  assign ram$206 = ram[206];
  assign ram$207 = ram[207];
  assign ram$208 = ram[208];
  assign ram$209 = ram[209];
  assign ram$210 = ram[210];
  assign ram$211 = ram[211];
  assign ram$212 = ram[212];
  assign ram$213 = ram[213];
  assign ram$214 = ram[214];
  assign ram$215 = ram[215];
  assign ram$216 = ram[216];
  assign ram$217 = ram[217];
  assign ram$218 = ram[218];
  assign ram$219 = ram[219];
  assign ram$220 = ram[220];
  assign ram$221 = ram[221];
  assign ram$222 = ram[222];
  assign ram$223 = ram[223];
  assign ram$224 = ram[224];
  assign ram$225 = ram[225];
  assign ram$226 = ram[226];
  assign ram$227 = ram[227];
  assign ram$228 = ram[228];
  assign ram$229 = ram[229];
  assign ram$230 = ram[230];
  assign ram$231 = ram[231];
  assign ram$232 = ram[232];
  assign ram$233 = ram[233];
  assign ram$234 = ram[234];
  assign ram$235 = ram[235];
  assign ram$236 = ram[236];
  assign ram$237 = ram[237];
  assign ram$238 = ram[238];
  assign ram$239 = ram[239];
  assign ram$240 = ram[240];
  assign ram$241 = ram[241];
  assign ram$242 = ram[242];
  assign ram$243 = ram[243];
  assign ram$244 = ram[244];
  assign ram$245 = ram[245];
  assign ram$246 = ram[246];
  assign ram$247 = ram[247];
  assign ram$248 = ram[248];
  assign ram$249 = ram[249];
  assign ram$250 = ram[250];
  assign ram$251 = ram[251];
  assign ram$252 = ram[252];
  assign ram$253 = ram[253];
  assign ram$254 = ram[254];
  assign ram$255 = ram[255];
  assign ram$256 = ram[256];
  assign ram$257 = ram[257];
  assign ram$258 = ram[258];
  assign ram$259 = ram[259];
  assign ram$260 = ram[260];
  assign ram$261 = ram[261];
  assign ram$262 = ram[262];
  assign ram$263 = ram[263];
  assign ram$264 = ram[264];
  assign ram$265 = ram[265];
  assign ram$266 = ram[266];
  assign ram$267 = ram[267];
  assign ram$268 = ram[268];
  assign ram$269 = ram[269];
  assign ram$270 = ram[270];
  assign ram$271 = ram[271];
  assign ram$272 = ram[272];
  assign ram$273 = ram[273];
  assign ram$274 = ram[274];
  assign ram$275 = ram[275];
  assign ram$276 = ram[276];
  assign ram$277 = ram[277];
  assign ram$278 = ram[278];
  assign ram$279 = ram[279];
  assign ram$280 = ram[280];
  assign ram$281 = ram[281];
  assign ram$282 = ram[282];
  assign ram$283 = ram[283];
  assign ram$284 = ram[284];
  assign ram$285 = ram[285];
  assign ram$286 = ram[286];
  assign ram$287 = ram[287];
  assign ram$288 = ram[288];
  assign ram$289 = ram[289];
  assign ram$290 = ram[290];
  assign ram$291 = ram[291];
  assign ram$292 = ram[292];
  assign ram$293 = ram[293];
  assign ram$294 = ram[294];
  assign ram$295 = ram[295];
  assign ram$296 = ram[296];
  assign ram$297 = ram[297];
  assign ram$298 = ram[298];
  assign ram$299 = ram[299];
  assign ram$300 = ram[300];
  assign ram$301 = ram[301];
  assign ram$302 = ram[302];
  assign ram$303 = ram[303];
  assign ram$304 = ram[304];
  assign ram$305 = ram[305];
  assign ram$306 = ram[306];
  assign ram$307 = ram[307];
  assign ram$308 = ram[308];
  assign ram$309 = ram[309];
  assign ram$310 = ram[310];
  assign ram$311 = ram[311];
  assign ram$312 = ram[312];
  assign ram$313 = ram[313];
  assign ram$314 = ram[314];
  assign ram$315 = ram[315];
  assign ram$316 = ram[316];
  assign ram$317 = ram[317];
  assign ram$318 = ram[318];
  assign ram$319 = ram[319];
  assign ram$320 = ram[320];
  assign ram$321 = ram[321];
  assign ram$322 = ram[322];
  assign ram$323 = ram[323];
  assign ram$324 = ram[324];
  assign ram$325 = ram[325];
  assign ram$326 = ram[326];
  assign ram$327 = ram[327];
  assign ram$328 = ram[328];
  assign ram$329 = ram[329];
  assign ram$330 = ram[330];
  assign ram$331 = ram[331];
  assign ram$332 = ram[332];
  assign ram$333 = ram[333];
  assign ram$334 = ram[334];
  assign ram$335 = ram[335];
  assign ram$336 = ram[336];
  assign ram$337 = ram[337];
  assign ram$338 = ram[338];
  assign ram$339 = ram[339];
  assign ram$340 = ram[340];
  assign ram$341 = ram[341];
  assign ram$342 = ram[342];
  assign ram$343 = ram[343];
  assign ram$344 = ram[344];
  assign ram$345 = ram[345];
  assign ram$346 = ram[346];
  assign ram$347 = ram[347];
  assign ram$348 = ram[348];
  assign ram$349 = ram[349];
  assign ram$350 = ram[350];
  assign ram$351 = ram[351];
  assign ram$352 = ram[352];
  assign ram$353 = ram[353];
  assign ram$354 = ram[354];
  assign ram$355 = ram[355];
  assign ram$356 = ram[356];
  assign ram$357 = ram[357];
  assign ram$358 = ram[358];
  assign ram$359 = ram[359];
  assign ram$360 = ram[360];
  assign ram$361 = ram[361];
  assign ram$362 = ram[362];
  assign ram$363 = ram[363];
  assign ram$364 = ram[364];
  assign ram$365 = ram[365];
  assign ram$366 = ram[366];
  assign ram$367 = ram[367];
  assign ram$368 = ram[368];
  assign ram$369 = ram[369];
  assign ram$370 = ram[370];
  assign ram$371 = ram[371];
  assign ram$372 = ram[372];
  assign ram$373 = ram[373];
  assign ram$374 = ram[374];
  assign ram$375 = ram[375];
  assign ram$376 = ram[376];
  assign ram$377 = ram[377];
  assign ram$378 = ram[378];
  assign ram$379 = ram[379];
  assign ram$380 = ram[380];
  assign ram$381 = ram[381];
  assign ram$382 = ram[382];
  assign ram$383 = ram[383];
  assign ram$384 = ram[384];
  assign ram$385 = ram[385];
  assign ram$386 = ram[386];
  assign ram$387 = ram[387];
  assign ram$388 = ram[388];
  assign ram$389 = ram[389];
  assign ram$390 = ram[390];
  assign ram$391 = ram[391];
  assign ram$392 = ram[392];
  assign ram$393 = ram[393];
  assign ram$394 = ram[394];
  assign ram$395 = ram[395];
  assign ram$396 = ram[396];
  assign ram$397 = ram[397];
  assign ram$398 = ram[398];
  assign ram$399 = ram[399];
  assign ram$400 = ram[400];
  assign ram$401 = ram[401];
  assign ram$402 = ram[402];
  assign ram$403 = ram[403];
  assign ram$404 = ram[404];
  assign ram$405 = ram[405];
  assign ram$406 = ram[406];
  assign ram$407 = ram[407];
  assign ram$408 = ram[408];
  assign ram$409 = ram[409];
  assign ram$410 = ram[410];
  assign ram$411 = ram[411];
  assign ram$412 = ram[412];
  assign ram$413 = ram[413];
  assign ram$414 = ram[414];
  assign ram$415 = ram[415];
  assign ram$416 = ram[416];
  assign ram$417 = ram[417];
  assign ram$418 = ram[418];
  assign ram$419 = ram[419];
  assign ram$420 = ram[420];
  assign ram$421 = ram[421];
  assign ram$422 = ram[422];
  assign ram$423 = ram[423];
  assign ram$424 = ram[424];
  assign ram$425 = ram[425];
  assign ram$426 = ram[426];
  assign ram$427 = ram[427];
  assign ram$428 = ram[428];
  assign ram$429 = ram[429];
  assign ram$430 = ram[430];
  assign ram$431 = ram[431];
  assign ram$432 = ram[432];
  assign ram$433 = ram[433];
  assign ram$434 = ram[434];
  assign ram$435 = ram[435];
  assign ram$436 = ram[436];
  assign ram$437 = ram[437];
  assign ram$438 = ram[438];
  assign ram$439 = ram[439];
  assign ram$440 = ram[440];
  assign ram$441 = ram[441];
  assign ram$442 = ram[442];
  assign ram$443 = ram[443];
  assign ram$444 = ram[444];
  assign ram$445 = ram[445];
  assign ram$446 = ram[446];
  assign ram$447 = ram[447];
  assign ram$448 = ram[448];
  assign ram$449 = ram[449];
  assign ram$450 = ram[450];
  assign ram$451 = ram[451];
  assign ram$452 = ram[452];
  assign ram$453 = ram[453];
  assign ram$454 = ram[454];
  assign ram$455 = ram[455];
  assign ram$456 = ram[456];
  assign ram$457 = ram[457];
  assign ram$458 = ram[458];
  assign ram$459 = ram[459];
  assign ram$460 = ram[460];
  assign ram$461 = ram[461];
  assign ram$462 = ram[462];
  assign ram$463 = ram[463];
  assign ram$464 = ram[464];
  assign ram$465 = ram[465];
  assign ram$466 = ram[466];
  assign ram$467 = ram[467];
  assign ram$468 = ram[468];
  assign ram$469 = ram[469];
  assign ram$470 = ram[470];
  assign ram$471 = ram[471];
  assign ram$472 = ram[472];
  assign ram$473 = ram[473];
  assign ram$474 = ram[474];
  assign ram$475 = ram[475];
  assign ram$476 = ram[476];
  assign ram$477 = ram[477];
  assign ram$478 = ram[478];
  assign ram$479 = ram[479];
  assign ram$480 = ram[480];
  assign ram$481 = ram[481];
  assign ram$482 = ram[482];
  assign ram$483 = ram[483];
  assign ram$484 = ram[484];
  assign ram$485 = ram[485];
  assign ram$486 = ram[486];
  assign ram$487 = ram[487];
  assign ram$488 = ram[488];
  assign ram$489 = ram[489];
  assign ram$490 = ram[490];
  assign ram$491 = ram[491];
  assign ram$492 = ram[492];
  assign ram$493 = ram[493];
  assign ram$494 = ram[494];
  assign ram$495 = ram[495];
  assign ram$496 = ram[496];
  assign ram$497 = ram[497];
  assign ram$498 = ram[498];
  assign ram$499 = ram[499];
  assign ram$500 = ram[500];
  assign ram$501 = ram[501];
  assign ram$502 = ram[502];
  assign ram$503 = ram[503];
  assign ram$504 = ram[504];
  assign ram$505 = ram[505];
  assign ram$506 = ram[506];
  assign ram$507 = ram[507];
  assign ram$508 = ram[508];
  assign ram$509 = ram[509];
  assign ram$510 = ram[510];
  assign ram$511 = ram[511];
  assign ram$512 = ram[512];
  assign ram$513 = ram[513];
  assign ram$514 = ram[514];
  assign ram$515 = ram[515];
  assign ram$516 = ram[516];
  assign ram$517 = ram[517];
  assign ram$518 = ram[518];
  assign ram$519 = ram[519];
  assign ram$520 = ram[520];
  assign ram$521 = ram[521];
  assign ram$522 = ram[522];
  assign ram$523 = ram[523];
  assign ram$524 = ram[524];
  assign ram$525 = ram[525];
  assign ram$526 = ram[526];
  assign ram$527 = ram[527];
  assign ram$528 = ram[528];
  assign ram$529 = ram[529];
  assign ram$530 = ram[530];
  assign ram$531 = ram[531];
  assign ram$532 = ram[532];
  assign ram$533 = ram[533];
  assign ram$534 = ram[534];
  assign ram$535 = ram[535];
  assign ram$536 = ram[536];
  assign ram$537 = ram[537];
  assign ram$538 = ram[538];
  assign ram$539 = ram[539];
  assign ram$540 = ram[540];
  assign ram$541 = ram[541];
  assign ram$542 = ram[542];
  assign ram$543 = ram[543];
  assign ram$544 = ram[544];
  assign ram$545 = ram[545];
  assign ram$546 = ram[546];
  assign ram$547 = ram[547];
  assign ram$548 = ram[548];
  assign ram$549 = ram[549];
  assign ram$550 = ram[550];
  assign ram$551 = ram[551];
  assign ram$552 = ram[552];
  assign ram$553 = ram[553];
  assign ram$554 = ram[554];
  assign ram$555 = ram[555];
  assign ram$556 = ram[556];
  assign ram$557 = ram[557];
  assign ram$558 = ram[558];
  assign ram$559 = ram[559];
  assign ram$560 = ram[560];
  assign ram$561 = ram[561];
  assign ram$562 = ram[562];
  assign ram$563 = ram[563];
  assign ram$564 = ram[564];
  assign ram$565 = ram[565];
  assign ram$566 = ram[566];
  assign ram$567 = ram[567];
  assign ram$568 = ram[568];
  assign ram$569 = ram[569];
  assign ram$570 = ram[570];
  assign ram$571 = ram[571];
  assign ram$572 = ram[572];
  assign ram$573 = ram[573];
  assign ram$574 = ram[574];
  assign ram$575 = ram[575];
  assign ram$576 = ram[576];
  assign ram$577 = ram[577];
  assign ram$578 = ram[578];
  assign ram$579 = ram[579];
  assign ram$580 = ram[580];
  assign ram$581 = ram[581];
  assign ram$582 = ram[582];
  assign ram$583 = ram[583];
  assign ram$584 = ram[584];
  assign ram$585 = ram[585];
  assign ram$586 = ram[586];
  assign ram$587 = ram[587];
  assign ram$588 = ram[588];
  assign ram$589 = ram[589];
  assign ram$590 = ram[590];
  assign ram$591 = ram[591];
  assign ram$592 = ram[592];
  assign ram$593 = ram[593];
  assign ram$594 = ram[594];
  assign ram$595 = ram[595];
  assign ram$596 = ram[596];
  assign ram$597 = ram[597];
  assign ram$598 = ram[598];
  assign ram$599 = ram[599];
  assign ram$600 = ram[600];
  assign ram$601 = ram[601];
  assign ram$602 = ram[602];
  assign ram$603 = ram[603];
  assign ram$604 = ram[604];
  assign ram$605 = ram[605];
  assign ram$606 = ram[606];
  assign ram$607 = ram[607];
  assign ram$608 = ram[608];
  assign ram$609 = ram[609];
  assign ram$610 = ram[610];
  assign ram$611 = ram[611];
  assign ram$612 = ram[612];
  assign ram$613 = ram[613];
  assign ram$614 = ram[614];
  assign ram$615 = ram[615];
  assign ram$616 = ram[616];
  assign ram$617 = ram[617];
  assign ram$618 = ram[618];
  assign ram$619 = ram[619];
  assign ram$620 = ram[620];
  assign ram$621 = ram[621];
  assign ram$622 = ram[622];
  assign ram$623 = ram[623];
  assign ram$624 = ram[624];
  assign ram$625 = ram[625];
  assign ram$626 = ram[626];
  assign ram$627 = ram[627];
  assign ram$628 = ram[628];
  assign ram$629 = ram[629];
  assign ram$630 = ram[630];
  assign ram$631 = ram[631];
  assign ram$632 = ram[632];
  assign ram$633 = ram[633];
  assign ram$634 = ram[634];
  assign ram$635 = ram[635];
  assign ram$636 = ram[636];
  assign ram$637 = ram[637];
  assign ram$638 = ram[638];
  assign ram$639 = ram[639];
  assign ram$640 = ram[640];
  assign ram$641 = ram[641];
  assign ram$642 = ram[642];
  assign ram$643 = ram[643];
  assign ram$644 = ram[644];
  assign ram$645 = ram[645];
  assign ram$646 = ram[646];
  assign ram$647 = ram[647];
  assign ram$648 = ram[648];
  assign ram$649 = ram[649];
  assign ram$650 = ram[650];
  assign ram$651 = ram[651];
  assign ram$652 = ram[652];
  assign ram$653 = ram[653];
  assign ram$654 = ram[654];
  assign ram$655 = ram[655];
  assign ram$656 = ram[656];
  assign ram$657 = ram[657];
  assign ram$658 = ram[658];
  assign ram$659 = ram[659];
  assign ram$660 = ram[660];
  assign ram$661 = ram[661];
  assign ram$662 = ram[662];
  assign ram$663 = ram[663];
  assign ram$664 = ram[664];
  assign ram$665 = ram[665];
  assign ram$666 = ram[666];
  assign ram$667 = ram[667];
  assign ram$668 = ram[668];
  assign ram$669 = ram[669];
  assign ram$670 = ram[670];
  assign ram$671 = ram[671];
  assign ram$672 = ram[672];
  assign ram$673 = ram[673];
  assign ram$674 = ram[674];
  assign ram$675 = ram[675];
  assign ram$676 = ram[676];
  assign ram$677 = ram[677];
  assign ram$678 = ram[678];
  assign ram$679 = ram[679];
  assign ram$680 = ram[680];
  assign ram$681 = ram[681];
  assign ram$682 = ram[682];
  assign ram$683 = ram[683];
  assign ram$684 = ram[684];
  assign ram$685 = ram[685];
  assign ram$686 = ram[686];
  assign ram$687 = ram[687];
  assign ram$688 = ram[688];
  assign ram$689 = ram[689];
  assign ram$690 = ram[690];
  assign ram$691 = ram[691];
  assign ram$692 = ram[692];
  assign ram$693 = ram[693];
  assign ram$694 = ram[694];
  assign ram$695 = ram[695];
  assign ram$696 = ram[696];
  assign ram$697 = ram[697];
  assign ram$698 = ram[698];
  assign ram$699 = ram[699];
  assign ram$700 = ram[700];
  assign ram$701 = ram[701];
  assign ram$702 = ram[702];
  assign ram$703 = ram[703];
  assign ram$704 = ram[704];
  assign ram$705 = ram[705];
  assign ram$706 = ram[706];
  assign ram$707 = ram[707];
  assign ram$708 = ram[708];
  assign ram$709 = ram[709];
  assign ram$710 = ram[710];
  assign ram$711 = ram[711];
  assign ram$712 = ram[712];
  assign ram$713 = ram[713];
  assign ram$714 = ram[714];
  assign ram$715 = ram[715];
  assign ram$716 = ram[716];
  assign ram$717 = ram[717];
  assign ram$718 = ram[718];
  assign ram$719 = ram[719];
  assign ram$720 = ram[720];
  assign ram$721 = ram[721];
  assign ram$722 = ram[722];
  assign ram$723 = ram[723];
  assign ram$724 = ram[724];
  assign ram$725 = ram[725];
  assign ram$726 = ram[726];
  assign ram$727 = ram[727];
  assign ram$728 = ram[728];
  assign ram$729 = ram[729];
  assign ram$730 = ram[730];
  assign ram$731 = ram[731];
  assign ram$732 = ram[732];
  assign ram$733 = ram[733];
  assign ram$734 = ram[734];
  assign ram$735 = ram[735];
  assign ram$736 = ram[736];
  assign ram$737 = ram[737];
  assign ram$738 = ram[738];
  assign ram$739 = ram[739];
  assign ram$740 = ram[740];
  assign ram$741 = ram[741];
  assign ram$742 = ram[742];
  assign ram$743 = ram[743];
  assign ram$744 = ram[744];
  assign ram$745 = ram[745];
  assign ram$746 = ram[746];
  assign ram$747 = ram[747];
  assign ram$748 = ram[748];
  assign ram$749 = ram[749];
  assign ram$750 = ram[750];
  assign ram$751 = ram[751];
  assign ram$752 = ram[752];
  assign ram$753 = ram[753];
  assign ram$754 = ram[754];
  assign ram$755 = ram[755];
  assign ram$756 = ram[756];
  assign ram$757 = ram[757];
  assign ram$758 = ram[758];
  assign ram$759 = ram[759];
  assign ram$760 = ram[760];
  assign ram$761 = ram[761];
  assign ram$762 = ram[762];
  assign ram$763 = ram[763];
  assign ram$764 = ram[764];
  assign ram$765 = ram[765];
  assign ram$766 = ram[766];
  assign ram$767 = ram[767];
  assign ram$768 = ram[768];
  assign ram$769 = ram[769];
  assign ram$770 = ram[770];
  assign ram$771 = ram[771];
  assign ram$772 = ram[772];
  assign ram$773 = ram[773];
  assign ram$774 = ram[774];
  assign ram$775 = ram[775];
  assign ram$776 = ram[776];
  assign ram$777 = ram[777];
  assign ram$778 = ram[778];
  assign ram$779 = ram[779];
  assign ram$780 = ram[780];
  assign ram$781 = ram[781];
  assign ram$782 = ram[782];
  assign ram$783 = ram[783];
  assign ram$784 = ram[784];
  assign ram$785 = ram[785];
  assign ram$786 = ram[786];
  assign ram$787 = ram[787];
  assign ram$788 = ram[788];
  assign ram$789 = ram[789];
  assign ram$790 = ram[790];
  assign ram$791 = ram[791];
  assign ram$792 = ram[792];
  assign ram$793 = ram[793];
  assign ram$794 = ram[794];
  assign ram$795 = ram[795];
  assign ram$796 = ram[796];
  assign ram$797 = ram[797];
  assign ram$798 = ram[798];
  assign ram$799 = ram[799];
  assign ram$800 = ram[800];
  assign ram$801 = ram[801];
  assign ram$802 = ram[802];
  assign ram$803 = ram[803];
  assign ram$804 = ram[804];
  assign ram$805 = ram[805];
  assign ram$806 = ram[806];
  assign ram$807 = ram[807];
  assign ram$808 = ram[808];
  assign ram$809 = ram[809];
  assign ram$810 = ram[810];
  assign ram$811 = ram[811];
  assign ram$812 = ram[812];
  assign ram$813 = ram[813];
  assign ram$814 = ram[814];
  assign ram$815 = ram[815];
  assign ram$816 = ram[816];
  assign ram$817 = ram[817];
  assign ram$818 = ram[818];
  assign ram$819 = ram[819];
  assign ram$820 = ram[820];
  assign ram$821 = ram[821];
  assign ram$822 = ram[822];
  assign ram$823 = ram[823];
  assign ram$824 = ram[824];
  assign ram$825 = ram[825];
  assign ram$826 = ram[826];
  assign ram$827 = ram[827];
  assign ram$828 = ram[828];
  assign ram$829 = ram[829];
  assign ram$830 = ram[830];
  assign ram$831 = ram[831];
  assign ram$832 = ram[832];
  assign ram$833 = ram[833];
  assign ram$834 = ram[834];
  assign ram$835 = ram[835];
  assign ram$836 = ram[836];
  assign ram$837 = ram[837];
  assign ram$838 = ram[838];
  assign ram$839 = ram[839];
  assign ram$840 = ram[840];
  assign ram$841 = ram[841];
  assign ram$842 = ram[842];
  assign ram$843 = ram[843];
  assign ram$844 = ram[844];
  assign ram$845 = ram[845];
  assign ram$846 = ram[846];
  assign ram$847 = ram[847];
  assign ram$848 = ram[848];
  assign ram$849 = ram[849];
  assign ram$850 = ram[850];
  assign ram$851 = ram[851];
  assign ram$852 = ram[852];
  assign ram$853 = ram[853];
  assign ram$854 = ram[854];
  assign ram$855 = ram[855];
  assign ram$856 = ram[856];
  assign ram$857 = ram[857];
  assign ram$858 = ram[858];
  assign ram$859 = ram[859];
  assign ram$860 = ram[860];
  assign ram$861 = ram[861];
  assign ram$862 = ram[862];
  assign ram$863 = ram[863];
  assign ram$864 = ram[864];
  assign ram$865 = ram[865];
  assign ram$866 = ram[866];
  assign ram$867 = ram[867];
  assign ram$868 = ram[868];
  assign ram$869 = ram[869];
  assign ram$870 = ram[870];
  assign ram$871 = ram[871];
  assign ram$872 = ram[872];
  assign ram$873 = ram[873];
  assign ram$874 = ram[874];
  assign ram$875 = ram[875];
  assign ram$876 = ram[876];
  assign ram$877 = ram[877];
  assign ram$878 = ram[878];
  assign ram$879 = ram[879];
  assign ram$880 = ram[880];
  assign ram$881 = ram[881];
  assign ram$882 = ram[882];
  assign ram$883 = ram[883];
  assign ram$884 = ram[884];
  assign ram$885 = ram[885];
  assign ram$886 = ram[886];
  assign ram$887 = ram[887];
  assign ram$888 = ram[888];
  assign ram$889 = ram[889];
  assign ram$890 = ram[890];
  assign ram$891 = ram[891];
  assign ram$892 = ram[892];
  assign ram$893 = ram[893];
  assign ram$894 = ram[894];
  assign ram$895 = ram[895];
  assign ram$896 = ram[896];
  assign ram$897 = ram[897];
  assign ram$898 = ram[898];
  assign ram$899 = ram[899];
  assign ram$900 = ram[900];
  assign ram$901 = ram[901];
  assign ram$902 = ram[902];
  assign ram$903 = ram[903];
  assign ram$904 = ram[904];
  assign ram$905 = ram[905];
  assign ram$906 = ram[906];
  assign ram$907 = ram[907];
  assign ram$908 = ram[908];
  assign ram$909 = ram[909];
  assign ram$910 = ram[910];
  assign ram$911 = ram[911];
  assign ram$912 = ram[912];
  assign ram$913 = ram[913];
  assign ram$914 = ram[914];
  assign ram$915 = ram[915];
  assign ram$916 = ram[916];
  assign ram$917 = ram[917];
  assign ram$918 = ram[918];
  assign ram$919 = ram[919];
  assign ram$920 = ram[920];
  assign ram$921 = ram[921];
  assign ram$922 = ram[922];
  assign ram$923 = ram[923];
  assign ram$924 = ram[924];
  assign ram$925 = ram[925];
  assign ram$926 = ram[926];
  assign ram$927 = ram[927];
  assign ram$928 = ram[928];
  assign ram$929 = ram[929];
  assign ram$930 = ram[930];
  assign ram$931 = ram[931];
  assign ram$932 = ram[932];
  assign ram$933 = ram[933];
  assign ram$934 = ram[934];
  assign ram$935 = ram[935];
  assign ram$936 = ram[936];
  assign ram$937 = ram[937];
  assign ram$938 = ram[938];
  assign ram$939 = ram[939];
  assign ram$940 = ram[940];
  assign ram$941 = ram[941];
  assign ram$942 = ram[942];
  assign ram$943 = ram[943];
  assign ram$944 = ram[944];
  assign ram$945 = ram[945];
  assign ram$946 = ram[946];
  assign ram$947 = ram[947];
  assign ram$948 = ram[948];
  assign ram$949 = ram[949];
  assign ram$950 = ram[950];
  assign ram$951 = ram[951];
  assign ram$952 = ram[952];
  assign ram$953 = ram[953];
  assign ram$954 = ram[954];
  assign ram$955 = ram[955];
  assign ram$956 = ram[956];
  assign ram$957 = ram[957];
  assign ram$958 = ram[958];
  assign ram$959 = ram[959];
  assign ram$960 = ram[960];
  assign ram$961 = ram[961];
  assign ram$962 = ram[962];
  assign ram$963 = ram[963];
  assign ram$964 = ram[964];
  assign ram$965 = ram[965];
  assign ram$966 = ram[966];
  assign ram$967 = ram[967];
  assign ram$968 = ram[968];
  assign ram$969 = ram[969];
  assign ram$970 = ram[970];
  assign ram$971 = ram[971];
  assign ram$972 = ram[972];
  assign ram$973 = ram[973];
  assign ram$974 = ram[974];
  assign ram$975 = ram[975];
  assign ram$976 = ram[976];
  assign ram$977 = ram[977];
  assign ram$978 = ram[978];
  assign ram$979 = ram[979];
  assign ram$980 = ram[980];
  assign ram$981 = ram[981];
  assign ram$982 = ram[982];
  assign ram$983 = ram[983];
  assign ram$984 = ram[984];
  assign ram$985 = ram[985];
  assign ram$986 = ram[986];
  assign ram$987 = ram[987];
  assign ram$988 = ram[988];
  assign ram$989 = ram[989];
  assign ram$990 = ram[990];
  assign ram$991 = ram[991];
  assign ram$992 = ram[992];
  assign ram$993 = ram[993];
  assign ram$994 = ram[994];
  assign ram$995 = ram[995];
  assign ram$996 = ram[996];
  assign ram$997 = ram[997];
  assign ram$998 = ram[998];
  assign ram$999 = ram[999];
  assign ram$1000 = ram[1000];
  assign ram$1001 = ram[1001];
  assign ram$1002 = ram[1002];
  assign ram$1003 = ram[1003];
  assign ram$1004 = ram[1004];
  assign ram$1005 = ram[1005];
  assign ram$1006 = ram[1006];
  assign ram$1007 = ram[1007];
  assign ram$1008 = ram[1008];
  assign ram$1009 = ram[1009];
  assign ram$1010 = ram[1010];
  assign ram$1011 = ram[1011];
  assign ram$1012 = ram[1012];
  assign ram$1013 = ram[1013];
  assign ram$1014 = ram[1014];
  assign ram$1015 = ram[1015];
  assign ram$1016 = ram[1016];
  assign ram$1017 = ram[1017];
  assign ram$1018 = ram[1018];
  assign ram$1019 = ram[1019];
  assign ram$1020 = ram[1020];
  assign ram$1021 = ram[1021];
  assign ram$1022 = ram[1022];
  assign ram$1023 = ram[1023];

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def port_a():
  //             if s.we_a:
  //                 s.ram[s.addr_a].next = s.data_a
  //                 s.q_a.next           = s.data_a
  //             else:
  //                 s.q_a.next = s.ram[s.addr_a]

  // logic for port_a()
  always @ (posedge clk) begin
    if (we_a) begin
      ram[addr_a] <= data_a;
      q_a <= data_a;
    end
    else begin
      q_a <= ram[addr_a];
    end
  //end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def port_b():
  //             if s.we_b:
  //                 s.ram[s.addr_b].next = s.data_b
  //                 s.q_b.next           = s.data_b
  //             else:
  //                 s.q_b.next = s.ram[s.addr_b]

  // logic for port_b()
  //always @ (posedge clk) begin
    if (we_b) begin
      ram[addr_b] <= data_b;
      q_b <= data_b;
    end
    else begin
      q_b <= ram[addr_b];
    end
  end


endmodule // ram_0x4915ea16bef085cd
`default_nettype wire

